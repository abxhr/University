// Code your design here
// Abshar Mohammed Aslam
// ID: 2019A7PS0233U

module NANDgate (A,B);
  input A;
  output B;
  
  nand (B,A,A);
endmodule