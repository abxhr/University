// Code your design here
// Abshar Mohammed Aslam
// ID: 2019A7PS0233U


module complement(x,y);
  input [7:0]x;
  output [7:0] y;
  assign y = ~x;
endmodule